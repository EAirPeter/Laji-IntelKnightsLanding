// dog auto generation
assign alu_data_res_ps3 = alu_data_res_ps2;
assign datamem_op_ps3 = datamem_op_ps2;
assign datamem_w_en_ps3 = datamem_w_en_ps2;
assign imm16_ps3 = imm16_ps2;
assign mux_regfile_data_w_ps3 = mux_regfile_data_w_ps2;
assign mux_regfile_req_w_ps3 = mux_regfile_req_w_ps2;
assign pc_4_ps3 = pc_4_ps2;
assign rd_ps3 = rd_ps2;
assign regfile_data_a_ps3 = regfile_data_a_ps2;
assign regfile_data_b_ps3 = regfile_data_b_ps2;
assign regfile_w_en_ps3 = regfile_w_en_ps2;
assign rt_ps3 = rt_ps2;
assign wtg_op_ps3 = wtg_op_ps2;
