// dog auto generation
assign inst_ps1 = inst_ps0;
assign pc_4_ps1 = pc_4_ps0;
