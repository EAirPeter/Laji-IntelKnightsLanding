`ifndef lajiintel_test_test_vh_
`define lajiintel_test_test_vh_

`include "../Auxiliary.vh"
`include "../Core.vh"

`define cp(x_)  #((x_) * 10)
`define ns(x_)  #(x_)
`define us(x_)  #((x_) * 1000)
`define ms(x_)  #((x_) * 1000_000)

`endif
