`undef GEN_F____
`undef GEN_FD___
`undef GEN_FDX__
`undef GEN_FDXM_
`undef GEN_FDXMW
`undef GEN_FDO__
`undef GEN_FDOM_
`undef GEN_FDOMW
`undef GEN__D___
`undef GEN__DX__
`undef GEN__DXM_
`undef GEN__DXMW
`undef GEN__DO__
`undef GEN__DOM_
`undef GEN__DOMW
`undef GEN___X__
`undef GEN___XM_
`undef GEN___XMW
`undef GEN____M_
`undef GEN____MW
`undef GEN_____W
