// dog auto generation
assign alu_op_ps2 = alu_op_ps1;
assign datamem_op_ps2 = datamem_op_ps1;
assign datamem_w_en_ps2 = datamem_w_en_ps1;
assign imm16_ps2 = imm16_ps1;
assign mux_alu_data_y_ps2 = mux_alu_data_y_ps1;
assign mux_regfile_data_w_ps2 = mux_regfile_data_w_ps1;
assign mux_regfile_req_w_ps2 = mux_regfile_req_w_ps1;
assign pc_4_ps2 = pc_4_ps1;
assign rd_ps2 = rd_ps1;
assign regfile_data_a_ps2 = regfile_data_a_ps1;
assign regfile_data_b_ps2 = regfile_data_b_ps1;
assign regfile_w_en_ps2 = regfile_w_en_ps1;
assign rt_ps2 = rt_ps1;
assign shamt_ps2 = shamt_ps1;
assign syscall_en_ps2 = syscall_en_ps1;
assign wtg_op_ps2 = wtg_op_ps1;
