// dog auto generation
assign alu_data_res_ps4 = alu_data_res_ps3;
assign datamem_data_ps4 = datamem_data_ps3;
assign mux_regfile_data_w_ps4 = mux_regfile_data_w_ps3;
assign mux_regfile_req_w_ps4 = mux_regfile_req_w_ps3;
assign pc_4_ps4 = pc_4_ps3;
assign rd_ps4 = rd_ps3;
assign regfile_w_en_ps4 = regfile_w_en_ps3;
assign rt_ps4 = rt_ps3;
